/*

//`resetall
//`timescale 1ns / 1ps
//`default_nettype none

/*
 * AXI4 2x2 interconnect (wrapper)
 */
module axi_interconnect_wrap_2x2 #
(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 32,
    parameter STRB_WIDTH = (DATA_WIDTH/8),
    parameter ID_WIDTH = 8,
    parameter M00_BASE_ADDR = 0,
    parameter M00_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M00_CONNECT_READ = 2'b11,
    parameter M00_CONNECT_WRITE = 2'b11,
    parameter M00_SECURE = 1'b0,
    parameter M01_BASE_ADDR = 0,
    parameter M01_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M01_CONNECT_READ = 2'b11,
    parameter M01_CONNECT_WRITE = 2'b11,
    parameter M01_SECURE = 1'b0
)
(
    input  wire                     clk,
    input  wire                     rst,

    /*
     * AXI slave interface
     */
    s00.axi_awid,
    s00.axi_awaddr,
    s00.axi_awlen,
    s00.axi_awsize,
    s00.axi_awburst,
    s00.axi_awlock,
    s00.axi_awcache,
    s00.axi_awprot,
    s00.axi_awqos,
    s00.axi_awuser,
    s00.axi_awvalid,
    s00.axi_awready,
    s00.axi_wdata,
    s00.axi_wstrb,
    s00.axi_wlast,
    s00.axi_wuser,
    s00.axi_wvalid,
    s00.axi_wready,
    s00.axi_bid,
    s00.axi_bresp,
    s00.axi_buser,
    s00.axi_bvalid,
    s00.axi_bready,
    s00.axi_arid,
    s00.axi_araddr,
    s00.axi_arlen,
    s00.axi_arsize,
    s00.axi_arburst,
    s00.axi_arlock,
    s00.axi_arcache,
    s00.axi_arprot,
    s00.axi_arqos,
    s00.axi_aruser,
    s00.axi_arvalid,
    s00.axi_arready,
    s00.axi_rid,
    s00.axi_rdata,
    s00.axi_rresp,
    s00.axi_rlast,
    s00.axi_ruser,
    s00.axi_rvalid,
    s00.axi_rready,

    s01.axi_awid,
    s01.axi_awaddr,
    s01.axi_awlen,
    s01.axi_awsize,
    s01.axi_awburst,
    s01.axi_awlock,
    s01.axi_awcache,
    s01.axi_awprot,
    s01.axi_awqos,
    s01.axi_awuser,
    s01.axi_awvalid,
    s01.axi_awready,
    s01.axi_wdata,
    s01.axi_wstrb,
    s01.axi_wlast,
    s01.axi_wuser,
    s01.axi_wvalid,
    s01.axi_wready,
    s01.axi_bid,
    s01.axi_bresp,
    s01.axi_buser,
    s01.axi_bvalid,
    s01.axi_bready,
    s01.axi_arid,
    s01.axi_araddr,
    s01.axi_arlen,
    s01.axi_arsize,
    s01.axi_arburst,
    s01.axi_arlock,
    s01.axi_arcache,
    s01.axi_arprot,
    s01.axi_arqos,
    s01.axi_aruser,
    s01.axi_arvalid,
    s01.axi_arready,
    s01.axi_rid,
    s01.axi_rdata,
    s01.axi_rresp,
    s01.axi_rlast,
    s01.axi_ruser,
    s01.axi_rvalid,
    s01.axi_rready,
                                     
    /*                                           
     * AXI master interface                      
     */                         
    m00.axi_awid,
    m00.axi_awaddr,
    m00.axi_awlen,
    m00.axi_awsize,
    m00.axi_awburst,
    m00.axi_awlock,
    m00.axi_awcache,
    m00.axi_awprot,
    m00.axi_awqos,
    m00.axi_awregion,
    m00.axi_awuser,
    m00.axi_awvalid,
    m00.axi_awready,
    m00.axi_wdata,
    m00.axi_wstrb,
    m00.axi_wlast,
    m00.axi_wuser,
    m00.axi_wvalid,
    m00.axi_wready,
    m00.axi_bid,
    m00.axi_bresp,
    m00.axi_buser,
    m00.axi_bvalid,
    m00.axi_bready,
    m00.axi_arid,
    m00.axi_araddr,
    m00.axi_arlen,
    m00.axi_arsize,
    m00.axi_arburst,
    m00.axi_arlock,
    m00.axi_arcache,
    m00.axi_arprot,
    m00.axi_arqos,
    m00.axi_arregion,
    m00.axi_aruser,
    m00.axi_arvalid,
    m00.axi_arready,
    m00.axi_rid,
    m00.axi_rdata,
    m00.axi_rresp,
    m00.axi_rlast,
    m00.axi_ruser,
    m00.axi_rvalid,
    m00.axi_rready,
                         
    m01.axi_awid,
    m01.axi_awaddr,
    m01.axi_awlen,
    m01.axi_awsize,
    m01.axi_awburst,
    m01.axi_awlock,
    m01.axi_awcache,
    m01.axi_awprot,
    m01.axi_awqos,
    m01.axi_awregion,
    m01.axi_awuser,
    m01.axi_awvalid,
    m01.axi_awready,
    m01.axi_wdata,
    m01.axi_wstrb,
    m01.axi_wlast,
    m01.axi_wuser,
    m01.axi_wvalid,
    m01.axi_wready,
    m01.axi_bid,
    m01.axi_bresp,
    m01.axi_buser,
    m01.axi_bvalid,
    m01.axi_bready,
    m01.axi_arid,
    m01.axi_araddr,
    m01.axi_arlen,
    m01.axi_arsize,
    m01.axi_arburst,
    m01.axi_arlock,
    m01.axi_arcache,
    m01.axi_arprot,
    m01.axi_arqos,
    m01.axi_arregion,
    m01.axi_aruser,
    m01.axi_arvalid,
    m01.axi_arready,
    m01.axi_rid,
    m01.axi_rdata,
    m01.axi_rresp,
    m01.axi_rlast,
    m01.axi_ruser,
    m01.axi_rvalid,
    m01.axi_rready
);

localparam S_COUNT = 2;
localparam M_COUNT = 2;

// parameter sizing helpers
function [ADDR_WIDTH*M_REGIONS-1:0] w_a_r(input [ADDR_WIDTH*M_REGIONS-1:0] val);
    w_a_r = val;
endfunction

function [32*M_REGIONS-1:0] w_32_r(input [32*M_REGIONS-1:0] val);
    w_32_r = val;
endfunction

function [S_COUNT-1:0] w_s(input [S_COUNT-1:0] val);
    w_s = val;
endfunction

function w_1(input val);
    w_1 = val;
endfunction

axi_interconnect #(
    .S_COUNT(S_COUNT),
    .M_COUNT(M_COUNT),
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(ADDR_WIDTH),
    .STRB_WIDTH(STRB_WIDTH),
    .ID_WIDTH(ID_WIDTH),
    .M_BASE_ADDR({ w_a_r(M01_BASE_ADDR), w_a_r(M00_BASE_ADDR) }),
    .M_ADDR_WIDTH({ w_32_r(M01_ADDR_WIDTH), w_32_r(M00_ADDR_WIDTH) }),
    .M_CONNECT_READ({ w_s(M01_CONNECT_READ), w_s(M00_CONNECT_READ) }),
    .M_CONNECT_WRITE({ w_s(M01_CONNECT_WRITE), w_s(M00_CONNECT_WRITE) }),
    .M_SECURE({ w_1(M01_SECURE), w_1(M00_SECURE) })
)
axi_interconnect_inst (
    .clk(clk),
    .rst(rst),
    .s_axi_awid({ s01.axi_awid, s00.axi_awid }),
    .s_axi_awaddr({ s01.axi_awaddr, s00.axi_awaddr }),
    .s_axi_awlen({ s01.axi_awlen, s00.axi_awlen }),
    .s_axi_awsize({ s01.axi_awsize, s00.axi_awsize }),
    .s_axi_awburst({ s01.axi_awburst, s00.axi_awburst }),
    .s_axi_awlock({ s01.axi_awlock, s00.axi_awlock }),
    .s_axi_awcache({ s01.axi_awcache, s00.axi_awcache }),
    .s_axi_awprot({ s01.axi_awprot, s00.axi_awprot }),
    .s_axi_awqos({ s01.axi_awqos, s00.axi_awqos }),
    .s_axi_awuser({ s01.axi_awuser, s00.axi_awuser }),
    .s_axi_awvalid({ s01.axi_awvalid, s00.axi_awvalid }),
    .s_axi_awready({ s01.axi_awready, s00.axi_awready }),
    .s_axi_wdata({ s01.axi_wdata, s00.axi_wdata }),
    .s_axi_wstrb({ s01.axi_wstrb, s00.axi_wstrb }),
    .s_axi_wlast({ s01.axi_wlast, s00.axi_wlast }),
    .s_axi_wuser({ s01.axi_wuser, s00.axi_wuser }),
    .s_axi_wvalid({ s01.axi_wvalid, s00.axi_wvalid }),
    .s_axi_wready({ s01.axi_wready, s00.axi_wready }),
    .s_axi_bid({ s01.axi_bid, s00.axi_bid }),
    .s_axi_bresp({ s01.axi_bresp, s00.axi_bresp }),
    .s_axi_buser({ s01.axi_buser, s00.axi_buser }),
    .s_axi_bvalid({ s01.axi_bvalid, s00.axi_bvalid }),
    .s_axi_bready({ s01.axi_bready, s00.axi_bready }),
    .s_axi_arid({ s01.axi_arid, s00.axi_arid }),
    .s_axi_araddr({ s01.axi_araddr, s00.axi_araddr }),
    .s_axi_arlen({ s01.axi_arlen, s00.axi_arlen }),
    .s_axi_arsize({ s01.axi_arsize, s00.axi_arsize }),
    .s_axi_arburst({ s01.axi_arburst, s00.axi_arburst }),
    .s_axi_arlock({ s01.axi_arlock, s00.axi_arlock }),
    .s_axi_arcache({ s01.axi_arcache, s00.axi_arcache }),
    .s_axi_arprot({ s01.axi_arprot, s00.axi_arprot }),
    .s_axi_arqos({ s01.axi_arqos, s00.axi_arqos }),
    .s_axi_aruser({ s01.axi_aruser, s00.axi_aruser }),
    .s_axi_arvalid({ s01.axi_arvalid, s00.axi_arvalid }),
    .s_axi_arready({ s01.axi_arready, s00.axi_arready }),
    .s_axi_rid({ s01.axi_rid, s00.axi_rid }),
    .s_axi_rdata({ s01.axi_rdata, s00.axi_rdata }),
    .s_axi_rresp({ s01.axi_rresp, s00.axi_rresp }),
    .s_axi_rlast({ s01.axi_rlast, s00.axi_rlast }),
    .s_axi_ruser({ s01.axi_ruser, s00.axi_ruser }),
    .s_axi_rvalid({ s01.axi_rvalid, s00.axi_rvalid }),
    .s_axi_rready({ s01.axi_rready, s00.axi_rready }),
    .m_axi_awid({ m01.axi_awid, m00.axi_awid }),
    .m_axi_awaddr({ m01.axi_awaddr, m00.axi_awaddr }),
    .m_axi_awlen({ m01.axi_awlen, m00.axi_awlen }),
    .m_axi_awsize({ m01.axi_awsize, m00.axi_awsize }),
    .m_axi_awburst({ m01.axi_awburst, m00.axi_awburst }),
    .m_axi_awlock({ m01.axi_awlock, m00.axi_awlock }),
    .m_axi_awcache({ m01.axi_awcache, m00.axi_awcache }),
    .m_axi_awprot({ m01.axi_awprot, m00.axi_awprot }),
    .m_axi_awqos({ m01.axi_awqos, m00.axi_awqos }),
    .m_axi_awregion({ m01.axi_awregion, m00.axi_awregion }),
    .m_axi_awuser({ m01.axi_awuser, m00.axi_awuser }),
    .m_axi_awvalid({ m01.axi_awvalid, m00.axi_awvalid }),
    .m_axi_awready({ m01.axi_awready, m00.axi_awready }),
    .m_axi_wdata({ m01.axi_wdata, m00.axi_wdata }),
    .m_axi_wstrb({ m01.axi_wstrb, m00.axi_wstrb }),
    .m_axi_wlast({ m01.axi_wlast, m00.axi_wlast }),
    .m_axi_wuser({ m01.axi_wuser, m00.axi_wuser }),
    .m_axi_wvalid({ m01.axi_wvalid, m00.axi_wvalid }),
    .m_axi_wready({ m01.axi_wready, m00.axi_wready }),
    .m_axi_bid({ m01.axi_bid, m00.axi_bid }),
    .m_axi_bresp({ m01.axi_bresp, m00.axi_bresp }),
    .m_axi_buser({ m01.axi_buser, m00.axi_buser }),
    .m_axi_bvalid({ m01.axi_bvalid, m00.axi_bvalid }),
    .m_axi_bready({ m01.axi_bready, m00.axi_bready }),
    .m_axi_arid({ m01.axi_arid, m00.axi_arid }),
    .m_axi_araddr({ m01.axi_araddr, m00.axi_araddr }),
    .m_axi_arlen({ m01.axi_arlen, m00.axi_arlen }),
    .m_axi_arsize({ m01.axi_arsize, m00.axi_arsize }),
    .m_axi_arburst({ m01.axi_arburst, m00.axi_arburst }),
    .m_axi_arlock({ m01.axi_arlock, m00.axi_arlock }),
    .m_axi_arcache({ m01.axi_arcache, m00.axi_arcache }),
    .m_axi_arprot({ m01.axi_arprot, m00.axi_arprot }),
    .m_axi_arqos({ m01.axi_arqos, m00.axi_arqos }),
    .m_axi_arregion({ m01.axi_arregion, m00.axi_arregion }),
    .m_axi_aruser({ m01.axi_aruser, m00.axi_aruser }),
    .m_axi_arvalid({ m01.axi_arvalid, m00.axi_arvalid }),
    .m_axi_arready({ m01.axi_arready, m00.axi_arready }),
    .m_axi_rid({ m01.axi_rid, m00.axi_rid }),
    .m_axi_rdata({ m01.axi_rdata, m00.axi_rdata }),
    .m_axi_rresp({ m01.axi_rresp, m00.axi_rresp }),
    .m_axi_rlast({ m01.axi_rlast, m00.axi_rlast }),
    .m_axi_ruser({ m01.axi_ruser, m00.axi_ruser }),
    .m_axi_rvalid({ m01.axi_rvalid, m00.axi_rvalid }),
    .m_axi_rready({ m01.axi_rready, m00.axi_rready })
);

endmodule

//`resetall
